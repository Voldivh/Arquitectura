//=======================================================
//  MODULE Definition
//=======================================================
module CSAI #(parameter DATAWIDTH_BUS=32)
(
	//////////// INPUTS //////////
	CLK, 
	RESET,
	ACK,
	CS,
	//////////// OUTPUTS //////////
	OUT
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
	input					 CLK;
	input					 RESET;
	input					 ACK;
	input			[10:0] CS;
	output reg	[10:0] OUT;
//=======================================================
//  REG/WIRE declarations
//=======================================================
//=======================================================
//  Structural coding
//=======================================================
// INPUT LOGIC: SEQUENTIAL
	always@(posedge CLK)
		begin 
			if(RESET == 1)
				OUT <= 0;
			else if(ACK==0)
				OUT = CS + 1;
			else
				OUT = CS;
		end
// INPUT LOGIC: COMBINATIONAL
//=======================================================
//  Outputs
//=======================================================
// OUTPUT LOGIC : COMBINATIONAL
endmodule
