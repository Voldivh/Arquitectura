
//=======================================================
//  MODULE Definition
//=======================================================
module MIR #(parameter DATAWIDTH_BUS_ADDRESS=11, DATAWIDTH_BUS_WORD=41)
(
	//////////// OUTPUTS //////////
	MIR_WORD,
	//////////// INPUTS //////////
	CLK,
	ADDRESS,
);
//=======================================================
//  PARAMETER declarations
//=======================================================

//=======================================================
//  PORT declarations
//=======================================================
	input		 CLK;
	input		[DATAWIDTH_BUS_ADDRESS-1:0] ADDRESS;
	
	output	[DATAWIDTH_BUS_WORD-1:0] MIR_WORD;
//=======================================================
//  REG/WIRE declarations
//=======================================================

	reg [DATAWIDTH_BUS_WORD-1:0] MIR_Register;
	reg [DATAWIDTH_BUS_WORD-1:0] MIR_Signal;

//=======================================================
//  Structural coding
//=======================================================
//INPUT LOGIC: COMBINATIONAL
	always@(ADDRESS)
		begin
			case (ADDRESS)

				11'd0    : MIR_Signal = 41'b00011000001100000111010010100000000000000; // Inicializar
				11'd1    : MIR_Signal = 41'b00000000000000000000000010111100000000000; // Decode
			
				// ADDCC
				11'd1600 : MIR_Signal = 41'b00000000000000000000000010110111001000010;//
				11'd1601 : MIR_Signal = 41'b00000010000001000000100001111011111111111; // 
				11'd1602 : MIR_Signal = 41'b00011100000000000101000110000000000000000; // 
				11'd1603 : MIR_Signal = 41'b00000010001010000000100001111011111111111; // 

				//be-ba
				11'd1088 : MIR_Signal = 41'b00000000000000000000000010111000000000010;// 
				11'd2	   : MIR_Signal = 41'b00011100000000000101000101000000000000000;//
				11'd3    : MIR_Signal = 41'b00010100000000000101000111100000000000000;// 
				11'd4    : MIR_Signal = 41'b00010100000000000101000111100000000000000;// 
				11'd5    : MIR_Signal = 41'b00011100000000000111000111100000000000000;// 
				11'd6	   : MIR_Signal = 41'b00011100000000000111000111100000000000000;//
				11'd7    : MIR_Signal = 41'b00011100000000000111000111100000000000000;//
				11'd8    : MIR_Signal = 41'b00011100001110000111000100010100000001100;// 
				11'd9    : MIR_Signal = 41'b00011100001110000111000100010100000001101;// 
				11'd10	: MIR_Signal = 41'b00011100001110000111000100001000000001100;//
				11'd11   : MIR_Signal = 41'b00000000000000000000000010111011111111111;// 
				11'd12   : MIR_Signal = 41'b00011000001010000110000100011000000000000;// 
				11'd13   : MIR_Signal = 41'b00011100001110000111000100010100000010000;// 
				11'd14   : MIR_Signal = 41'b00000000000000000000000010110000000001100;//
				11'd15   : MIR_Signal = 41'b00000000000000000000000010111011111111111;// 
				11'd16   : MIR_Signal = 41'b00000000000000000000000010110100000010011;// 
				11'd17   : MIR_Signal = 41'b00000000000000000000000010100100000001100;//
				11'd18   : MIR_Signal = 41'b00000000000000000000000010111011111111111;// 
				11'd19   : MIR_Signal = 41'b00000000000000000000000010101100000001100;// 
				11'd20   : MIR_Signal = 41'b00000000000000000000000010111011111111111;// 
				
				// SUBCC
				11'd1584 : MIR_Signal = 41'b00011100000000000101000110010111000110010;//
				11'd1585 : MIR_Signal = 41'b00000000000001000101000100000000000000000;// 
				11'd1586 : MIR_Signal = 41'b00010100000000000101000011100000000000000;//
				11'd1587 : MIR_Signal = 41'b00010100000000000101000110111011001000011;// 
				
				11'd2047 : MIR_Signal = 41'b00011000000000000110000111011000000000000;
				
				default: MIR_Signal = MIR_Register; // 
			endcase
		end
		
//STATE REGISTER: SEQUENTIAL
	always @(posedge CLK)
	begin
			MIR_Register <= MIR_Signal;
	end
//=======================================================
//  Outputs
//=======================================================
// OUTPUT LOGIC : COMBINATIONAL
assign MIR_WORD = MIR_Register;

endmodule